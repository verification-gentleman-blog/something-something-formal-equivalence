// Copyright 2020 Tudor Timisescu (verificationgentleman.com)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


module equivalence_tb(
    input bit PCLK,
    input bit PRESETn,
    input struct {
      bit PSEL;
      bit PENABLE;
      bit PWRITE;
      bit [31:0] PWDATA;
      bit [3:0] PSTRB;
    } sigs[2]);

  for (genvar i = 0; i < 2; i++) begin: duts
    dummy dut(
        .PCLK(PCLK),
        .PRESETn(PRESETn),
        .PSEL(sigs[i].PSEL),
        .PENABLE(sigs[i].PENABLE),
        .PWRITE(sigs[i].PWRITE),
        .PWDATA(sigs[i].PWDATA),
        .PSTRB(sigs[i].PSTRB));
  end

endmodule
